module xilix_bram_tdp
#(  // Parameters
    parameter         BRAM_SIZE             = "36Kb",        // Target BRAM: "18Kb" or "36Kb"
    parameter integer PORT_A_OUT_REG        = 1,             // Optional port A output register (0 or 1)
    parameter integer PORT_B_OUT_REG        = 1,             // Optional port B output register (0 or 1)
    parameter integer INIT_A                = 36'd0,         // Initial values on port A output port
    parameter integer INIT_B                = 36'd0,         // Initial values on port B output port
    parameter         INIT_FILE             = "NONE",                  
    parameter integer READ_WIDTH_A          = 16,            // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
    parameter integer READ_WIDTH_B          = 16,            // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
    parameter         SIM_COLLISION_CHK     = "ALL",         // Collision check enable "ALL", "WARNING_ONLY", // "GENERATE_X_ONLY" or "NONE"
    parameter integer SRVAL_A               = 36'd0,         // Set/Reset value for port A output
    parameter integer SRVAL_B               = 36'd0,         // Set/Reset value for port B output
    parameter         WRITE_MODE_A          = "WRITE_FIRST", // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
    parameter         WRITE_MODE_B          = "WRITE_FIRST", // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
    parameter         WRITE_WIDTH_A         = 16,            // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
    parameter         WRITE_WIDTH_B         = 16             // Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
)(  //Ports                                                  
    output wire [ READ_WIDTH_A    -1 : 0 ]  DOA,             // Output port-A data, width defined by READ_WIDTH_A parameter
    output wire [ READ_WIDTH_B    -1 : 0 ]  DOB,             // Output port-B data, width defined by READ_WIDTH_B parameter
    input  wire [ ADDRA_WIDTH     -1 : 0 ]  ADDRA,           // Input port-A address, width defined by Port A depth
    input  wire [ ADDRB_WIDTH     -1 : 0 ]  ADDRB,           // Input port-B address, width defined by Port B depth
    input  wire                             CLKA,            // 1-bit input port-A clock
    input  wire                             CLKB,            // 1-bit input port-B clock
    input  wire [ WRITE_WIDTH_A   -1 : 0 ]  DIA,             // Input port-A data, width defined by WRITE_WIDTH_A parameter
    input  wire [ WRITE_WIDTH_B   -1 : 0 ]  DIB,             // Input port-B data, width defined by WRITE_WIDTH_B parameter
    input  wire                             ENA,             // 1-bit input port-A enable
    input  wire                             ENB,             // 1-bit input port-B enable
    input  wire                             REGCEA,          // 1-bit input port-A output register enable
    input  wire                             REGCEB,          // 1-bit input port-B output register enable
    input  wire                             RSTA,            // 1-bit input port-A reset
    input  wire                             RSTB,            // 1-bit input port-B reset
    input  wire [ WEA_WIDTH       -1 : 0 ]  WEA,             // Input port-A write enable, width defined by Port A depth
    input  wire [ WEB_WIDTH       -1 : 0 ]  WEB              // Input port-B write enable, width defined by Port B depth
);

localparam least_width_A =  (READ_WIDTH_A <= WRITE_WIDTH_A) ? READ_WIDTH_A : WRITE_WIDTH_A;
localparam least_width_B =  (READ_WIDTH_B <= WRITE_WIDTH_B) ? READ_WIDTH_B : WRITE_WIDTH_B;
localparam ADDRA_WIDTH   =  (BRAM_SIZE == "9Kb") ? ( (least_width_A == 1) ? 13 : (least_width_A == 2) ? 12 : (least_width_A > 2 && least_width_A <= 4) ? 11 : (least_width_A > 4 && least_width_A <= 9) ? 10 : (least_width_A > 9 && least_width_A <= 18) ? 9 : 13 ) : (BRAM_SIZE == "18Kb") ? ( (least_width_A == 1) ? 14 : (least_width_A == 2) ? 13 : (least_width_A > 2 && least_width_A <= 4) ? 12 : (least_width_A > 4 && least_width_A <= 9) ? 11 : (least_width_A > 9 && least_width_A <= 18) ? 10 : (least_width_A > 18 && least_width_A < 36) ? 9 : 14 ) : (BRAM_SIZE == "36Kb") ? ( (least_width_A == 1) ? 15 : (least_width_A == 2) ? 14 : (least_width_A > 2 && least_width_A <= 4) ? 13 : (least_width_A > 4 && least_width_A <= 9) ? 12 : (least_width_A > 9 && least_width_A <= 18) ? 11 : (least_width_A > 18 && least_width_A <= 36) ? 10 : 15 ) : 15;
localparam ADDRB_WIDTH   = (BRAM_SIZE == "9Kb") ? ( (least_width_B == 1) ? 13 : (least_width_B == 2) ? 12 : (least_width_B > 2 && least_width_B <= 4) ? 11 : (least_width_B > 4 && least_width_B <= 9) ? 10 : (least_width_B > 9 && least_width_B <= 18) ? 9 : 13 ) : (BRAM_SIZE == "18Kb") ? ( (least_width_B == 1) ? 14 : (least_width_B == 2) ? 13 : (least_width_B > 2 && least_width_B <= 4) ? 12 : (least_width_B > 4 && least_width_B <= 9) ? 11 : (least_width_B > 9 && least_width_B <= 18) ? 10 : (least_width_B > 18 && least_width_B <= 36 ) ? 9 : 14 ) : (BRAM_SIZE == "36Kb") ? ( (least_width_B == 1) ? 15 : (least_width_B == 2) ? 14 : (least_width_B > 2 && least_width_B <= 4) ? 13 : (least_width_B > 4 && least_width_B <= 9) ? 12 : (least_width_B > 9 && least_width_B <= 18) ? 11 : (least_width_B > 18 && least_width_B <= 36) ? 10 : 15 ) : 15;


localparam WEA_WIDTH = (WRITE_WIDTH_A <= 9) ? 1 : (WRITE_WIDTH_A > 9 && WRITE_WIDTH_A <= 18) ? 2 : (WRITE_WIDTH_A > 18 && WRITE_WIDTH_A <= 36) ? 4 : (BRAM_SIZE == "18Kb") ? 2 : 4;
localparam WEB_WIDTH = (WRITE_WIDTH_B <= 9) ? 1 : (WRITE_WIDTH_B > 9 && WRITE_WIDTH_B <= 18) ? 2 : (WRITE_WIDTH_B > 18 && WRITE_WIDTH_B <= 36) ? 4 : (BRAM_SIZE == "18Kb") ? 2 : 4;

// ******************************************************************
// MACRO: TRUE DUAL PORT BRAM
// ******************************************************************
BRAM_TDP_MACRO #(
    .BRAM_SIZE              ( BRAM_SIZE         ), 
    .DEVICE                 ( "7SERIES"         ), 
    .DOA_REG                ( PORT_A_OUT_REG    ), 
    .DOB_REG                ( PORT_B_OUT_REG    ), 
    .INIT_A                 ( INIT_A            ), 
    .INIT_B                 ( INIT_B            ), 
    .INIT_FILE              ( INIT_FILE         ),
    .READ_WIDTH_A           ( READ_WIDTH_A      ), 
    .READ_WIDTH_B           ( READ_WIDTH_B      ), 
    .SIM_COLLISION_CHECK    ( SIM_COLLISION_CHK ), 
    .SRVAL_A                ( SRVAL_A           ), 
    .SRVAL_B                ( SRVAL_B           ), 
    .WRITE_MODE_A           ( WRITE_MODE_A      ), 
    .WRITE_MODE_B           ( WRITE_MODE_B      ), 
    .WRITE_WIDTH_A          ( WRITE_WIDTH_A     ), 
    .WRITE_WIDTH_B          ( WRITE_WIDTH_B     )  
) BRAM_TDP_MACRO_inst (
    .DOA                    ( DOA               ), 
    .DOB                    ( DOB               ), 
    .ADDRA                  ( ADDRA             ), 
    .ADDRB                  ( ADDRB             ), 
    .CLKA                   ( CLKA              ), 
    .CLKB                   ( CLKB              ), 
    .DIA                    ( DIA               ), 
    .DIB                    ( DIB               ), 
    .ENA                    ( ENA               ), 
    .ENB                    ( ENB               ), 
    .REGCEA                 ( REGCEA            ), 
    .REGCEB                 ( REGCEB            ), 
    .RSTA                   ( RSTA              ), 
    .RSTB                   ( RSTB              ), 
    .WEA                    ( WEA               ), 
    .WEB                    ( WEB               )  
);

endmodule



    //// .INIT_00                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_01                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_02                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_03                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_04                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_05                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_06                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_07                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_08                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_09                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_0A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_0B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_0C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_0D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_0E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_0F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_10                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_11                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_12                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_13                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_14                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_15                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_16                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_17                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_18                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_19                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_1A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_1B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_1C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_1D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_1E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_1F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_20                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_21                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_22                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_23                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_24                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_25                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_26                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_27                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_28                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_29                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_2A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_2B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_2C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_2D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_2E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_2F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_30                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_31                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_32                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_33                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_34                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_35                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_36                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_37                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_38                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_39                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_3A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_3B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_3C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_3D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_3E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_3F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// // The next set of INIT_xx are valid when configured as 36Kb
    //// .INIT_40                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_41                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_42                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_43                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_44                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_45                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_46                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_47                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_48                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_49                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_4A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_4B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_4C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_4D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_4E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_4F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_50                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_51                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_52                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_53                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_54                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_55                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_56                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_57                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_58                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_59                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_5A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_5B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_5C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_5D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_5E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_5F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_60                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_61                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_62                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_63                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_64                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_65                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_66                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_67                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_68                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_69                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_6A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_6B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_6C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_6D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_6E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_6F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_70                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_71                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_72                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_73                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_74                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_75                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_76                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_77                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_78                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_79                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_7A                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_7B                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_7C                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_7D                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_7E                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INIT_7F                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),

    //// // The next set of INITP_xx are for the parity bits
    //// .INIT_FF                ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_00               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_01               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_02               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_03               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_04               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_05               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_06               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_07               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// // The next set of INITP_xx are valid when configured as 36Kb
    //// .INITP_08               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_09               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_0A               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_0B               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_0C               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_0D               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_0E               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    //// .INITP_0F               ( 256'h0000000000000000000000000000000000000000000000000000000000000000 )

