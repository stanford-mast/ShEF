001000001000000001100000101111010000000000000110000000000001000000001100000000000000000000000000000000000001101100000000100000000000000000000000000001001100000001000000000100
000100001000000000100000001111010000000000000010000000000001000000000100000000000000000000000000010011000000101100000000000000000000000000000000000011000100000001000000000100
001000001000000000100000000000000100000001111101000000000000000000100000000000000000000000001100100000000000000000000000000000000000000000000000000011111000000000000000000000
001000001000000000100000000000000100000000000010100000000000000000100000000000000000000000000111110100000000000000000000000000000000000000000000000000000100000000000000000000
