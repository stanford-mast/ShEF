0000000001000000000000011100000000000000000000001100000000000000000000000000011000000000000000000000000000000000010011
0000000001000000000010010100000000000000000000000001000000000000000000000000000010000000000000000000000000000000110001
0100000001000000010101110110000000000000000000011111100000000000000000000000111111000000000000000000000000000000000000
0100000001000010010000111001000000000000000000000001000000000000000000000000000010000000000000000000000000000000000000
