000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100
000000000001000000000000000000000000000000000000000000000000001111110000000000000000000000000000000100000000000000000000000000011100000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000010100000000000000000000000000000000010000000000000000000000000000010100000000000000000000000000000101
000000000001000000000000011100000000000000000000000000000000001111110000000000000000000000000001010000000000000000000000000000001100000000000000000000000000000011000000000000000000000001010000000000000000000000000000000000110010000000000000000000000000000101000000000000000000000000000000010100000000000000000000000000000101
000100000001000000000010010100000000000000000000000000000000001111110000000000000000000000000011001000000000000000000000000000000100000000000000000000000000000001000000000000000000111111110000000000000000000000000000000111110100000000000000000000000000000000010000000000000000000000110010000000000000000000000000000000000001
000100000001000000010101110110000000000000000000000000000000001111110000000000000000000000011111010000000000000000000000000000000001000000000000000000000000000000010000000000001101010100001111000000000000000000000000000000001010000000000000000000000000000000010000000000000000000000011111010000000000000000000000000000000001
