module stream_read_tb;

  reg clk;
  reg rst_n;
  reg  [31:0]  tb_req_addr;
  reg  [8:0]   tb_req_burst_count;
  reg          tb_req_val;
  wire         tb_req_rdy;

  wire [63:0] s_axi_rdata;
  wire s_axi_rvalid;
  reg  s_axi_rready;

  wire [15:0]  m_axi_arid;
  wire [63:0]  m_axi_araddr;
  wire [7:0]   m_axi_arlen;
  wire [2:0]   m_axi_arsize;
  wire [1:0]   m_axi_arburst;
  wire [1:0]   m_axi_arlock;
  wire [3:0]   m_axi_arcache;
  wire [2:0]   m_axi_arprot;
  wire [3:0]   m_axi_arqos;
  wire [3:0]   m_axi_arregion;
  wire         m_axi_arvalid;
  wire         m_axi_arready;
  wire [15:0]  m_axi_rid;
  wire [511:0] m_axi_rdata;
  wire [1:0]   m_axi_rresp;
  wire         m_axi_rlast;
  wire         m_axi_rvalid;
  wire         m_axi_rready;

  // ******************************************************************
  // Clock generation
  // ******************************************************************
  always begin : clk_gen
    #5;
    clk = !clk;
  end

  // ******************************************************************
  // DUT
  // ******************************************************************
  //
  stream_read dut(
    .clk(clk),
    .rst_n(rst_n),
    .req_addr(tb_req_addr),
    .req_burst_count(tb_req_burst_count),
    .req_val(tb_req_val),
    .req_rdy(tb_req_rdy),
    .s_axi_rid(), //SET TO 0
    .s_axi_rdata(s_axi_rdata),
    .s_axi_rresp(), //ALWAYS SUCCESS
    .s_axi_rlast(), //IGNORE FOR NOW
    .s_axi_rvalid(s_axi_rvalid),
    .s_axi_rready(s_axi_rready),
    .m_axi_arid    (m_axi_arid    ),
    .m_axi_araddr  (m_axi_araddr  ),
    .m_axi_arlen   (m_axi_arlen   ),
    .m_axi_arsize  (m_axi_arsize  ),
    .m_axi_arburst (m_axi_arburst ),
    .m_axi_arlock  (m_axi_arlock  ),
    .m_axi_arcache (m_axi_arcache ),
    .m_axi_arprot  (m_axi_arprot  ),
    .m_axi_arqos   (m_axi_arqos   ),
    .m_axi_arregion(m_axi_arregion),
    .m_axi_arvalid (m_axi_arvalid ),
    .m_axi_arready (m_axi_arready ),
    .m_axi_rid     (m_axi_rid     ),
    .m_axi_rdata   (m_axi_rdata   ),
    .m_axi_rresp   (m_axi_rresp   ),
    .m_axi_rlast   (m_axi_rlast   ),
    .m_axi_rvalid  (m_axi_rvalid  ),
    .m_axi_rready  (m_axi_rready  )
  );


  axi_driver axi_driver_inst(
    .clk(clk),
    .reset(~rst_n),
    .M_AXI_AWID       (),
    .M_AXI_AWADDR     (),
    .M_AXI_AWLEN      (),
    .M_AXI_AWSIZE     (),
    .M_AXI_AWBURST    (),
    .M_AXI_AWLOCK     (),
    .M_AXI_AWCACHE    (),
    .M_AXI_AWPROT     (),
    .M_AXI_AWQOS      (),
    .M_AXI_AWVALID    (),
    .M_AXI_AWREADY    (),
    .M_AXI_WID        (),
    .M_AXI_WDATA      (),
    .M_AXI_WSTRB      (),
    .M_AXI_WLAST      (),
    .M_AXI_WVALID     (),
    .M_AXI_WREADY     (),
    .M_AXI_BID        (),
    .M_AXI_BRESP      (),
    .M_AXI_BVALID     (),
    .M_AXI_BREADY     (),
    .M_AXI_ARID       (m_axi_arid    ),
    .M_AXI_ARADDR     (m_axi_araddr  ),
    .M_AXI_ARLEN      (m_axi_arlen   ),
    .M_AXI_ARSIZE     (m_axi_arsize  ),
    .M_AXI_ARBURST    (m_axi_arburst ),
    .M_AXI_ARLOCK     (m_axi_arlock  ),
    .M_AXI_ARCACHE    (m_axi_arcache ),
    .M_AXI_ARPROT     (m_axi_arprot  ),
    .M_AXI_ARQOS      (m_axi_arqos   ),
    .M_AXI_ARVALID    (m_axi_arvalid ),
    .M_AXI_ARREADY    (m_axi_arready ),
    .M_AXI_RID        (m_axi_rid     ),
    .M_AXI_RDATA      (m_axi_rdata   ),
    .M_AXI_RRESP      (m_axi_rresp   ),
    .M_AXI_RLAST      (m_axi_rlast   ),
    .M_AXI_RVALID     (m_axi_rvalid  ),
    .M_AXI_RREADY     (m_axi_rready  )
  );

  // ******************************************************************
  // Tasks
  // ******************************************************************
  task init_sim;
    begin
      clk = 1'b0;
      rst_n = 1'b1;

      tb_req_addr = 0;
      tb_req_burst_count = 0;
      tb_req_val = 0;
      s_axi_rready = 0;
    end
  endtask

  task reset_dut;
    begin
      $display("**** Toggling reset **** ");
      rst_n = 1'b0;

      #20;
      rst_n = 1'b1;
      @(posedge clk);
      $display("Reset done at %0t",$time);
    end
  endtask

  task read_burst;
    input [31:0] addr;
    input [7:0] burst_count;
    input [63:0] expected;
    reg [63:0] data;
    begin
      $display("Reading %d bursts from address %x", burst_count, addr);

      @(posedge clk);
      //Make the request
      tb_req_val = 1'b1;
      tb_req_addr = addr;
      tb_req_burst_count = burst_count;
      wait(tb_req_rdy);
      @(negedge clk);
      @(negedge clk);
      tb_req_val = 1'b0;

      @(posedge clk);

      for(int i = 0; i < burst_count; i++) begin
        s_axi_rready = 1'b1;
        #1;
        wait(s_axi_rvalid);
        @(negedge clk);
        data = s_axi_rdata;
        @(posedge clk);
        s_axi_rready = 1'b0;
        $display("      Read data: %x, expected %x", data, expected);
        if(data != expected) begin
          $display("     ERROR");
          $finish;
        end
      end
      $display("    OK");
    end
  endtask

  initial begin
    $display("***************************************");
    $display ("Testing read stream");
    $display("***************************************");
    init_sim();
    reset_dut();
    
    #20;

    read_burst(32'h0, 8'h1, 64'h0);
    //Read burst of longer than 1
    read_burst(32'h0, 8'h4, 64'h0);
    //Read burst that goes over one line
    read_burst(32'h0, 8'h9, 64'h0);
    
    //Read burst that is unaligned
    read_burst(32'h0000_0008, 8'h1, 64'h0); //still in line 0, should be muxed
    read_burst(32'h0000_0040, 8'h1, 64'h0); //index into ram line 1
    //Unaligned, multiple lines
    read_burst(32'h0000_0830, 8'd17, 64'h0); //over 3 lines. 2 bursts from first line, 8 from second, 7 from last
    
    //Evict
    read_burst(32'h0000_1000, 8'd1, 64'h0000_1000);
    read_burst(32'h0000_1ff8, 8'd1, 64'h0000_1000);
    
    read_burst(32'h0f00_3ff8, 8'd1, 64'h0f00_3000); //Evict with unaligned addr
    read_burst(32'h0f00_3030, 8'd15, 64'h0f00_3000);
    read_burst(32'h0f00_3000, 8'd1, 64'h0f00_3000);
    read_burst(32'h0000_0008, 8'h1, 64'h0);
    

    #100;
    $finish;
  end

endmodule
